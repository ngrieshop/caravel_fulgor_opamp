magic
tech sky130A
magscale 1 2
timestamp 1608352248
<< nwell >>
rect -5252 1004 -4822 1124
rect -5252 694 -4826 1004
<< pwell >>
rect -5252 504 -4822 546
rect -5252 192 -4826 504
rect -5252 188 -5242 192
rect -5182 188 -4826 192
<< psubdiff >>
rect -5252 240 -5188 294
rect -4884 240 -4822 294
<< nsubdiff >>
rect -5214 974 -5188 1028
rect -4884 974 -4860 1028
<< psubdiffcont >>
rect -5188 240 -4884 294
<< nsubdiffcont >>
rect -5188 974 -4884 1028
<< poly >>
rect -5048 650 -5018 931
rect -5180 634 -5018 650
rect -5180 594 -5164 634
rect -5084 594 -5018 634
rect -5180 576 -5018 594
rect -5048 351 -5018 576
<< polycont >>
rect -5164 594 -5084 634
<< locali >>
rect -5252 974 -5188 1028
rect -4884 974 -4822 1028
rect -5180 634 -5066 650
rect -5180 594 -5164 634
rect -5084 594 -5066 634
rect -5180 576 -5066 594
rect -5252 240 -5188 294
rect -4884 240 -4822 294
<< viali >>
rect -5164 594 -5084 634
<< metal1 >>
rect -5252 944 -4822 1056
rect -5096 826 -5062 944
rect -5006 650 -4971 838
rect -5252 634 -5066 650
rect -5252 594 -5164 634
rect -5084 594 -5066 634
rect -5252 576 -5066 594
rect -5006 576 -4822 650
rect -5132 408 -5122 484
rect -5070 408 -5060 484
rect -5006 373 -4971 576
rect -5252 228 -4822 332
<< via1 >>
rect -5122 408 -5070 484
<< metal2 >>
rect -5122 484 -5070 494
rect -5252 408 -5122 482
rect -5070 408 -4822 482
rect -5252 396 -4822 408
use sky130_fd_pr__pfet_01v8_35M7SK  sky130_fd_pr__pfet_01v8_35M7SK_0
timestamp 1608326616
transform 1 0 -5033 0 1 822
box -211 -128 211 188
use sky130_fd_pr__nfet_01v8_PUCP6T  inv_nfet
timestamp 1608326735
transform 1 0 -5033 0 1 443
box -211 -255 211 77
<< end >>
