**.subckt ring_vco
x1 10 out_ring o1 9 not
V1 vss GND DC{Vss} 
V2 vdd vss DC{Vdd} 
x2 10 o1 o2 9 not
x3 10 o2 o3 9 not
x4 10 o3 o4 9 not
x5 10 o4 o5 9 not
x6 10 o5 o6 9 not
XM1 out_ring o6 9 9 sky130_fd_pr__nfet_01v8 W=1.2 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XM2 out_ring o6 10 10 sky130_fd_pr__pfet_01v8 W=1.2 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XM3 out out_ring vss vss sky130_fd_pr__nfet_01v8 W=0.6 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XM4 out out_ring vdd vdd sky130_fd_pr__pfet_01v8 W=1.05 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XM5 10 5 vdd vdd sky130_fd_pr__pfet_01v8 W=1.2 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XM6 9 in vss vss sky130_fd_pr__nfet_01v8 W=1.2 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XM7 5 5 vdd vdd sky130_fd_pr__pfet_01v8 W=1.2 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XM8 5 in vss vss sky130_fd_pr__nfet_01v8 W=1.2 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
V3 in vss DC{Vin} 
**** begin user architecture code




* Circuit Parameters
.param vdd  = 1.8
.param vss  = 0.0
.param vin  = 0.3
.param iref = 200u
.options TEMP = 65.0

* Include Models
.lib ~/skywater_pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/sky130.lib TT

* OP Parameters & Singals to save
.save all  @M.X1.XM1.msky130_fd_pr__nfet_01v8[id] @M.X1.XM1.msky130_fd_pr__nfet_01v8[vth]
+ @M.X1.XM1.msky130_fd_pr__nfet_01v8[vgs] @M.X1.XM1.msky130_fd_pr__nfet_01v8[vds] @M.X1.XM1.msky130_fd_pr__nfet_01v8[vdsat]
+ @M.X1.XM1.msky130_fd_pr__nfet_01v8[gm] @M.X1.XM1.msky130_fd_pr__nfet_01v8[gds]  @M.X1.XM2.msky130_fd_pr__pfet_01v8[id]
+ @M.X1.XM2.msky130_fd_pr__pfet_01v8[vth] @M.X1.XM2.msky130_fd_pr__pfet_01v8[vgs] @M.X1.XM2.msky130_fd_pr__pfet_01v8[vds]
+ @M.X1.XM2.msky130_fd_pr__pfet_01v8[vdsat] @M.X1.XM2.msky130_fd_pr__pfet_01v8[gm] @M.X1.XM2.msky130_fd_pr__pfet_01v8[gds]

*Simulations
.control
  *reset
  tran 0.1n 0.5u
  stop when time = 0.1u
  alterparam vin = 1.8
  resume
  setplot tran1
  plot v(out)
  *write ~/caravel_fulgor_opamp/xschem/sim_results/opamp_closeloop_tran1.raw


  *dc V3 0 1.8 0.01
  *setplot dc1
  *plot v(out1) v(out2) v(out3) v(in)

  reset
  op
  setplot op1

.endc

.end


**** end user architecture code
**.ends

* expanding   symbol:  /home/dhernando/caravel_fulgor_opamp/xschem/ring_vco/not.sym # of pins=4

.subckt not  vdd in out vss
*.ipin vdd
*.ipin in
*.ipin vss
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8 W=0.42 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 W=0.42 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
.ends

.GLOBAL GND
.end
