magic
tech sky130A
magscale 1 2
timestamp 1608255475
<< error_s >>
rect -660 4266 -658 4449
rect -670 4263 -658 4266
rect -675 4251 -658 4263
rect -1220 3794 -1203 3806
rect -1220 3791 -1208 3794
rect -1220 3581 -1218 3791
rect -1220 3578 -1208 3581
rect -1220 3566 -1203 3578
<< nwell >>
rect -5124 5190 -146 5532
rect -764 4923 -438 4926
rect -1025 4454 -438 4923
rect -1444 4440 -438 4454
rect -1444 4032 -603 4440
<< pwell >>
rect -1443 3778 -433 4011
rect -1446 3356 -433 3778
rect -5124 2464 -134 2800
<< psubdiff >>
rect -4962 2652 -4902 2692
rect -3534 2652 -3488 2692
rect -4964 2556 -4904 2596
rect -3536 2556 -3490 2596
<< nsubdiff >>
rect -4908 5400 -4866 5440
rect -3574 5400 -3540 5440
rect -4912 5304 -4870 5344
rect -3578 5304 -3544 5344
<< psubdiffcont >>
rect -4902 2652 -3534 2692
rect -4904 2556 -3536 2596
<< nsubdiffcont >>
rect -4866 5400 -3574 5440
rect -4870 5304 -3578 5344
<< poly >>
rect -1248 3557 -1218 4431
rect -660 3722 -630 4449
<< locali >>
rect -4908 5400 -4866 5440
rect -3574 5400 -3540 5440
rect -4912 5304 -4870 5344
rect -3578 5304 -3544 5344
rect -4962 2652 -4902 2692
rect -3534 2652 -3488 2692
rect -4964 2556 -4904 2596
rect -3536 2556 -3490 2596
<< metal1 >>
rect -5122 5198 -144 5516
rect -4874 5051 -4832 5198
rect -4804 5082 -4794 5142
rect -4734 5082 -4724 5142
rect -4874 4888 -4790 5051
rect -3768 5046 -3726 5198
rect -3698 5088 -3688 5148
rect -3628 5088 -3618 5148
rect -4726 5040 -4470 5046
rect -4874 4886 -4832 4888
rect -4896 3112 -4822 3114
rect -4898 2932 -4822 3112
rect -4736 3109 -4470 5040
rect -3768 4849 -3698 5046
rect -3636 4526 -3499 5046
rect -4256 4306 -1718 4526
rect -4256 4280 -1722 4306
rect -4256 4172 -4036 4280
rect -3636 4240 -3566 4280
rect -1834 4172 -1722 4280
rect -4767 2937 -4470 3109
rect -3770 2956 -3696 3138
rect -4736 2935 -4470 2937
rect -4898 2804 -4862 2932
rect -4834 2848 -4824 2902
rect -4764 2848 -4754 2902
rect -3768 2804 -3732 2956
rect -3640 2950 -3608 3532
rect -3702 2844 -3692 2898
rect -3632 2844 -3622 2898
rect -5118 2642 -136 2804
rect -5118 2624 -132 2642
rect -5114 2462 -132 2624
<< via1 >>
rect -4794 5082 -4734 5142
rect -3688 5088 -3628 5148
rect -4824 2848 -4764 2902
rect -3692 2844 -3632 2898
<< metal2 >>
rect -4794 5148 -4734 5152
rect -3688 5148 -3628 5158
rect -4802 5142 -3688 5148
rect -4802 5090 -4794 5142
rect -4734 5090 -3688 5142
rect -4794 5072 -4734 5082
rect -3688 5078 -3628 5088
rect -4824 2910 -4764 2912
rect -4836 2902 -3632 2910
rect -4836 2848 -4824 2902
rect -4764 2898 -3632 2902
rect -4764 2848 -3692 2898
rect -4824 2838 -4764 2848
rect -3692 2834 -3632 2844
use via_li_m1  via_li_m1_1
array 0 19 72 0 0 74
timestamp 1607692587
transform 1 0 -4942 0 1 2536
box 4 0 76 74
use inverter  inverter_1
array 0 4 502 0 0 1206
timestamp 1608252737
transform 1 0 990 0 1 3228
box -5287 266 -4718 1124
use via_li_m1  via_li_m1_0
array 0 19 72 0 0 74
timestamp 1607692587
transform 1 0 -4942 0 1 2636
box 4 0 76 74
use sky130_fd_pr__nfet_01v8_YK3456  sky130_fd_pr__nfet_01v8_YK3456_0
timestamp 1608249442
transform -1 0 -4795 0 -1 3024
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_ZE46K8  sky130_fd_pr__nfet_01v8_ZE46K8_0
timestamp 1608249480
transform -1 0 -3669 0 -1 3045
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_3D5K6R  sky130_fd_pr__pfet_01v8_3D5K6R_0
timestamp 1608253231
transform 1 0 -3667 0 1 4954
box -211 -324 211 324
use sky130_fd_pr__pfet_01v8_35M7SK  sky130_fd_pr__pfet_01v8_35M7SK_0
timestamp 1608253040
transform -1 0 -4765 0 1 4961
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_373K6R  sky130_fd_pr__pfet_01v8_373K6R_0
timestamp 1608255150
transform 1 0 -643 0 1 4359
box -211 -327 211 327
use sky130_fd_pr__nfet_01v8_9TXQ83  sky130_fd_pr__nfet_01v8_9TXQ83_1
timestamp 1608229483
transform 1 0 -645 0 1 3648
box -211 -264 211 264
use sky130_fd_pr__nfet_01v8_R7545W  sky130_fd_pr__nfet_01v8_R7545W_0
timestamp 1608229183
transform 1 0 -1235 0 1 3686
box -211 -330 211 330
use sky130_fd_pr__pfet_01v8_3FZUWK  sky130_fd_pr__pfet_01v8_3FZUWK_0
timestamp 1608254796
transform 1 0 -1233 0 1 4468
box -211 -436 211 459
use via_li_m1  via_li_m1_3
array 0 19 72 0 0 74
timestamp 1607692587
transform 1 0 -4914 0 1 5286
box 4 0 76 74
use via_li_m1  via_li_m1_2
array 0 19 72 0 0 74
timestamp 1607692587
transform 1 0 -4906 0 1 5386
box 4 0 76 74
<< end >>
