magic
tech sky130A
magscale 1 2
timestamp 1608334096
<< nwell >>
rect -704 1454 2933 1455
rect -704 1114 2935 1454
rect -704 996 549 1114
rect 673 996 2935 1114
rect -704 665 2935 996
rect -704 662 2933 665
<< pwell >>
rect -692 619 2939 620
rect -692 -9 2941 619
rect -509 -10 2941 -9
<< metal1 >>
rect -601 1175 2846 1360
rect 558 1012 568 1101
rect 635 1012 645 1101
rect 1731 1004 1741 1110
rect 1841 1004 1851 1110
rect -704 612 -694 698
rect -626 612 -616 698
rect 2275 695 2285 724
rect -17 603 -7 687
rect 84 603 94 687
rect 538 616 860 667
rect 908 627 1242 690
rect 1713 632 2027 683
rect 2090 632 2285 695
rect 2275 616 2285 632
rect 2386 695 2396 724
rect 2386 632 2454 695
rect 2386 616 2396 632
rect 544 298 554 374
rect 634 298 644 374
rect 1734 306 1744 382
rect 1797 306 1807 382
rect -580 53 2876 242
<< via1 >>
rect 568 1012 635 1101
rect 1741 1004 1841 1110
rect -694 612 -626 698
rect -7 603 84 687
rect 2285 616 2386 724
rect 554 298 634 374
rect 1744 306 1797 382
<< metal2 >>
rect -165 1100 -80 1110
rect -165 999 -80 1009
rect 568 1101 635 1111
rect 568 1002 635 1012
rect 1741 1110 1841 1120
rect -697 890 -621 900
rect -697 768 -621 778
rect -692 708 -631 768
rect -694 698 -626 708
rect -694 602 -626 612
rect -692 537 -631 602
rect -700 527 -621 537
rect -700 437 -621 447
rect -159 379 -89 999
rect 568 881 632 1002
rect 1741 994 1841 1004
rect 555 871 647 881
rect 555 774 647 784
rect 568 761 632 774
rect 2285 724 2386 734
rect -22 687 91 698
rect -22 603 -7 687
rect 84 603 91 687
rect 2285 606 2386 616
rect 2846 696 2956 713
rect 2846 621 2862 696
rect 2939 621 2956 696
rect -22 592 91 603
rect 1732 533 1806 543
rect 2293 526 2377 606
rect 2846 596 2956 621
rect 1732 453 1806 463
rect 2283 516 2395 526
rect -166 369 -61 379
rect 554 374 634 384
rect 554 288 634 298
rect 1743 382 1798 453
rect 2283 399 2395 409
rect 1743 306 1744 382
rect 1797 306 1798 382
rect 1743 296 1798 306
rect -166 268 -61 278
<< via2 >>
rect -165 1009 -80 1100
rect 1741 1004 1841 1110
rect -697 778 -621 890
rect -700 447 -621 527
rect 555 784 647 871
rect -7 603 84 687
rect 2862 621 2939 696
rect 1732 463 1806 533
rect -166 278 -61 369
rect 554 298 634 374
rect 2283 409 2395 516
<< metal3 >>
rect 1731 1110 1851 1115
rect -175 1100 -70 1105
rect -175 1009 -165 1100
rect -80 1093 -70 1100
rect 1731 1093 1741 1110
rect -80 1014 1741 1093
rect -80 1009 -70 1014
rect -175 1004 -70 1009
rect 1731 1004 1741 1014
rect 1841 1004 1851 1110
rect 1731 999 1851 1004
rect -707 890 -611 895
rect -707 778 -697 890
rect -621 885 -611 890
rect -621 876 641 885
rect -621 871 657 876
rect -621 785 555 871
rect -621 778 -611 785
rect 545 784 555 785
rect 647 784 657 871
rect 545 779 657 784
rect -707 773 -611 778
rect -40 709 96 716
rect -40 696 2960 709
rect -40 687 2862 696
rect -40 603 -7 687
rect 84 621 2862 687
rect 2939 621 2960 696
rect 84 604 2960 621
rect 84 603 96 604
rect -40 584 96 603
rect 1722 533 1816 538
rect -710 527 -611 532
rect -710 447 -700 527
rect -621 523 -611 527
rect 1722 523 1732 533
rect -621 463 1732 523
rect 1806 523 1816 533
rect 1806 463 1817 523
rect 2273 517 2405 521
rect -621 452 1817 463
rect 2272 516 3151 517
rect -621 447 -611 452
rect -710 442 -611 447
rect 2272 409 2283 516
rect 2395 409 3151 516
rect 2272 407 3151 409
rect 2273 404 2405 407
rect -161 374 649 381
rect -176 369 554 374
rect -176 278 -166 369
rect -61 298 554 369
rect 634 298 649 374
rect -61 287 649 298
rect -61 278 -51 287
rect -176 273 -51 278
use inverter_fd  inverter_fd_0
timestamp 1608331766
transform 1 0 -456 0 1 -20
box 456 20 1060 1458
use trans_gate  trans_gate_0
timestamp 1608331766
transform 1 0 738 0 1 710
box -157 -701 436 733
use inverter_fd  inverter_fd_1
timestamp 1608331766
transform 1 0 712 0 1 -8
box 456 20 1060 1458
use trans_gate  trans_gate_1
timestamp 1608331766
transform 1 0 1913 0 1 718
box -157 -701 436 733
use inverter_fd  inverter_fd_2
timestamp 1608331766
transform 1 0 1876 0 1 -3
box 456 20 1060 1458
use inverter_fd  inverter_fd_3
timestamp 1608331766
transform 1 0 -1147 0 1 -17
box 456 20 1060 1458
<< labels >>
rlabel metal3 2395 407 3151 517 1 out
rlabel via1 -694 612 -626 698 1 in
rlabel metal1 -580 53 2876 242 1 vss
rlabel nwell -601 1175 2847 1360 1 vdd
<< end >>
