magic
tech sky130A
magscale 1 2
timestamp 1608340837
<< nwell >>
rect 3563 672 3809 1469
rect 3572 -1405 3818 -608
<< pwell >>
rect 3626 75 3793 614
rect 3626 67 3650 75
rect 3588 -550 3755 55
<< metal1 >>
rect -186 1368 675 1370
rect -278 1185 675 1368
rect 2942 1190 4485 1375
rect -278 -1126 -97 1185
rect 6464 233 7624 257
rect 64 -203 7624 233
rect 7437 -224 7624 -203
rect -278 -1160 2469 -1126
rect 2915 -1160 4402 -1126
rect -278 -1654 5306 -1160
rect -278 -1676 2469 -1654
rect -218 -1679 2469 -1676
rect -222 -2258 -212 -2144
rect -56 -2157 -46 -2144
rect -56 -2173 1869 -2157
rect -56 -2236 2008 -2173
rect -56 -2251 1869 -2236
rect -56 -2258 -46 -2251
rect 7437 -2612 7626 -224
rect 4717 -2801 7626 -2612
<< via1 >>
rect -212 -2258 -56 -2144
<< metal2 >>
rect 6 722 96 732
rect 6 588 96 598
rect 7359 539 7473 549
rect 7332 401 7359 493
rect 7332 391 7473 401
rect -208 -338 -88 -328
rect -208 -498 -88 -488
rect -204 -692 -96 -498
rect -203 -2134 -96 -692
rect 7332 -717 7465 391
rect -212 -2144 -56 -2134
rect -212 -2268 -56 -2258
rect -203 -2272 -96 -2268
<< via2 >>
rect 6 598 96 722
rect 7359 401 7473 539
rect -208 -488 -88 -338
<< metal3 >>
rect -10 732 116 926
rect -296 722 116 732
rect -296 610 6 722
rect -10 598 6 610
rect 96 598 116 722
rect -10 442 116 598
rect 7349 539 7483 544
rect 7349 401 7359 539
rect 7473 401 7483 539
rect 7349 396 7483 401
rect -218 -338 -78 -333
rect -218 -488 -208 -338
rect -88 -488 -78 -338
rect -218 -493 -78 -488
rect 5415 -2447 7363 -2337
use freq_div  freq_div_4
timestamp 1608334096
transform 1 0 2484 0 1 -2854
box -710 -10 3151 1455
use freq_div  freq_div_0
timestamp 1608334096
transform 1 0 710 0 1 10
box -710 -10 3151 1455
use freq_div  freq_div_1
timestamp 1608334096
transform 1 0 4426 0 1 15
box -710 -10 3151 1455
use freq_div  freq_div_3
timestamp 1608334096
transform -1 0 6671 0 -1 54
box -710 -10 3151 1455
use freq_div  freq_div_2
timestamp 1608334096
transform -1 0 2955 0 -1 49
box -710 -10 3151 1455
<< labels >>
rlabel metal3 -296 610 116 732 1 in
rlabel space 4879 -2447 7363 -2337 1 out
rlabel space 1904 -2801 7626 -2612 1 vss
rlabel space 2942 1190 7273 1375 1 vdd
<< end >>
