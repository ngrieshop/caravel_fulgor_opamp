magic
tech sky130A
magscale 1 2
timestamp 1608348248
<< nwell >>
rect -4208 9978 7720 11293
<< metal1 >>
rect 5922 12160 6111 12370
rect 5508 12087 8474 12160
rect 5331 11745 8474 12087
rect 5508 11700 8474 11745
rect -4208 10010 7689 10710
rect -4144 9957 7593 10010
rect -4281 8521 -4271 8612
rect -4133 8521 -4123 8612
rect 8124 7463 8466 11700
rect 7366 7121 8466 7463
<< via1 >>
rect -4271 8521 -4133 8612
<< metal2 >>
rect 5575 14223 5805 15861
rect -4257 11354 -4151 11364
rect -4257 11205 -4151 11215
rect -4251 8622 -4157 11205
rect -4271 8612 -4133 8622
rect -4271 8511 -4133 8521
rect -4251 8487 -4157 8511
rect -4332 7988 -4252 7998
rect -4332 7894 -4252 7904
rect 4885 7568 5059 7627
rect 2693 7512 7358 7568
rect 4885 6001 5059 7512
<< via2 >>
rect -4257 11215 -4151 11354
rect -4332 7904 -4252 7988
<< metal3 >>
rect -4267 11354 -4141 11359
rect -4267 11347 -4257 11354
rect -4551 11225 -4257 11347
rect -4267 11215 -4257 11225
rect -4151 11347 -4141 11354
rect -4151 11225 -1526 11347
rect -4151 11215 -4141 11225
rect -4267 11210 -4141 11215
rect -4502 7988 -4234 7998
rect -4502 7904 -4332 7988
rect -4252 7904 -4234 7988
rect -4502 7900 -4234 7904
rect -4342 7899 -4242 7900
use ring_vco  ring_vco_0
timestamp 1608340973
transform -1 0 2594 0 1 4659
box -5124 2462 6897 5532
use divx32  divx32_0
timestamp 1608345554
transform 1 0 -1515 0 -1 11957
box -296 -3279 7626 1470
<< labels >>
rlabel metal3 -4551 11225 -4429 11347 1 vco_out
rlabel metal3 -4502 7900 -4332 7998 1 enable
rlabel metal2 4885 6001 5059 7627 1 in
rlabel metal2 5575 15631 5805 15861 1 out_div
rlabel space -1793 9857 5758 10767 1 vdd
rlabel space -1733 13083 5028 13636 1 vdd
rlabel space -4204 7123 7718 7459 1 vss
rlabel space -1451 11724 8474 12160 1 vss
rlabel space 389 14569 3835 15168 1 vss
<< end >>
