magic
tech sky130A
magscale 1 2
timestamp 1608329555
<< error_s >>
rect -5124 5190 -4300 5403
rect -3685 3922 -3578 4160
rect -3116 3922 -3009 4160
rect -2547 3922 -2440 4160
rect -1978 3922 -1871 4160
rect -1409 3922 -1302 4160
rect -840 3922 -733 4160
rect -271 3922 -164 4160
rect 298 3922 405 4160
rect 867 3922 974 4160
rect 1436 3922 1543 4160
rect 2005 3922 2112 4160
rect 2574 3922 2681 4160
rect 3143 3922 3250 4160
rect 3712 3922 3819 4160
rect 4281 3922 4388 4160
rect 4850 3922 4957 4160
rect 5419 3922 5526 4160
rect 5988 3922 6095 4160
rect 6557 3922 6664 4160
rect 7126 3922 7233 4160
<< nwell >>
rect 8339 5532 9230 5539
rect -5124 5192 9230 5532
rect -5124 5190 8274 5192
rect 7802 4352 8106 4888
rect 8339 4870 8442 4884
rect 8135 4352 8400 4870
rect -4314 4350 7650 4352
rect -4256 4160 7650 4350
rect 7700 4160 8400 4352
rect 8054 3926 8400 4160
rect 8732 3924 9228 5192
<< pwell >>
rect 8006 3903 8400 3908
rect 7999 3670 8400 3903
rect 7996 3248 8400 3670
rect 8006 3228 8400 3248
rect 7928 3220 8400 3228
rect 8602 3220 9258 3906
rect 8132 2800 9260 3220
rect -5124 2464 9268 2800
<< psubdiff >>
rect 8150 3154 8210 3190
rect 9074 3154 9160 3190
rect 8154 3052 8214 3088
rect 9078 3052 9164 3088
rect 8156 2958 8216 2994
rect 9080 2958 9166 2994
rect 8156 2846 8216 2882
rect 9080 2846 9166 2882
rect -4962 2652 -4902 2692
rect -3534 2652 -3488 2692
rect -3072 2666 -3012 2706
rect -1644 2666 -1598 2706
rect -440 2676 -380 2716
rect 988 2676 1034 2716
rect 2298 2666 2358 2706
rect 3726 2666 3772 2706
rect 7708 2694 7768 2734
rect 9136 2694 9182 2734
rect 4998 2638 5058 2678
rect 6426 2638 6472 2678
rect -4964 2556 -4904 2596
rect -3536 2556 -3490 2596
rect -3074 2570 -3014 2610
rect -1646 2570 -1600 2610
rect -442 2580 -382 2620
rect 986 2580 1032 2620
rect 2296 2570 2356 2610
rect 3724 2570 3770 2610
rect 7706 2598 7766 2638
rect 9134 2598 9180 2638
rect 4996 2542 5056 2582
rect 6424 2542 6470 2582
<< nsubdiff >>
rect -4908 5400 -4866 5440
rect -3574 5400 -3540 5440
rect -2724 5404 -2682 5444
rect -1390 5404 -1356 5444
rect -92 5394 -50 5434
rect 1242 5394 1276 5434
rect 2266 5422 2308 5462
rect 3600 5422 3634 5462
rect 4890 5394 4932 5434
rect 6224 5394 6258 5434
rect 7238 5422 7280 5462
rect 8572 5422 8606 5462
rect -4912 5304 -4870 5344
rect -3578 5304 -3544 5344
rect -2728 5308 -2686 5348
rect -1394 5308 -1360 5348
rect -96 5298 -54 5338
rect 1238 5298 1272 5338
rect 2262 5326 2304 5366
rect 3596 5326 3630 5366
rect 4886 5298 4928 5338
rect 6220 5298 6254 5338
rect 7234 5326 7276 5366
rect 8568 5326 8602 5366
rect 7908 4700 7982 4740
rect 7908 4452 7982 4516
rect 7714 4222 7778 4296
rect 7962 4222 8002 4296
<< psubdiffcont >>
rect 8210 3154 9074 3190
rect 8214 3052 9078 3088
rect 8216 2958 9080 2994
rect 8216 2846 9080 2882
rect -4902 2652 -3534 2692
rect -3012 2666 -1644 2706
rect -380 2676 988 2716
rect 2358 2666 3726 2706
rect 7768 2694 9136 2734
rect 5058 2638 6426 2678
rect -4904 2556 -3536 2596
rect -3014 2570 -1646 2610
rect -382 2580 986 2620
rect 2356 2570 3724 2610
rect 7766 2598 9134 2638
rect 5056 2542 6424 2582
<< nsubdiffcont >>
rect -4866 5400 -3574 5440
rect -2682 5404 -1390 5444
rect -50 5394 1242 5434
rect 2308 5422 3600 5462
rect 4932 5394 6224 5434
rect 7280 5422 8572 5462
rect -4870 5304 -3578 5344
rect -2686 5308 -1394 5348
rect -54 5298 1238 5338
rect 2304 5326 3596 5366
rect 4928 5298 6220 5338
rect 7276 5326 8568 5366
rect 7908 4516 7982 4700
rect 7778 4222 7962 4296
<< poly >>
rect 8216 3920 8246 4699
rect 8659 3936 8689 3953
rect 7594 3886 8246 3920
rect 8216 3371 8246 3886
rect 8624 3920 8689 3936
rect 9008 3920 9038 4403
rect 8624 3886 9038 3920
rect 8624 3870 8689 3886
rect 8659 3857 8689 3870
rect 9008 3485 9038 3886
<< locali >>
rect -4908 5400 -4866 5440
rect -3574 5400 -3540 5440
rect -2724 5410 -2710 5444
rect -1380 5410 -1342 5444
rect -1308 5410 -1278 5444
rect -2724 5404 -2682 5410
rect -1390 5404 -1356 5410
rect -92 5400 -78 5434
rect 1252 5400 1290 5434
rect 1324 5400 1354 5434
rect 2266 5428 2280 5462
rect 3610 5428 3648 5462
rect 3682 5428 3712 5462
rect 2266 5422 2308 5428
rect 3600 5422 3634 5428
rect 4890 5400 4904 5434
rect 6234 5400 6272 5434
rect 6306 5400 6336 5434
rect 7238 5428 7252 5462
rect 8582 5428 8620 5462
rect 8654 5428 8684 5462
rect 7238 5422 7280 5428
rect 8572 5422 8606 5428
rect -92 5394 -50 5400
rect 1242 5394 1276 5400
rect 4890 5394 4932 5400
rect 6224 5394 6258 5400
rect 2262 5362 2304 5366
rect 3596 5362 3630 5366
rect 7234 5362 7276 5366
rect 8568 5362 8602 5366
rect -2728 5344 -2686 5348
rect -1394 5344 -1360 5348
rect -4912 5304 -4870 5344
rect -3578 5304 -3544 5344
rect -2728 5310 -2718 5344
rect -1388 5310 -1350 5344
rect -1316 5310 -1286 5344
rect -96 5334 -54 5338
rect 1238 5334 1272 5338
rect -2728 5308 -2686 5310
rect -1394 5308 -1360 5310
rect -96 5300 -86 5334
rect 1244 5300 1282 5334
rect 1316 5300 1346 5334
rect 2262 5328 2272 5362
rect 3602 5328 3640 5362
rect 3674 5328 3704 5362
rect 4886 5334 4928 5338
rect 6220 5334 6254 5338
rect 2262 5326 2304 5328
rect 3596 5326 3630 5328
rect 4886 5300 4896 5334
rect 6226 5300 6264 5334
rect 6298 5300 6328 5334
rect 7234 5328 7244 5362
rect 8574 5328 8612 5362
rect 8646 5328 8676 5362
rect 7234 5326 7276 5328
rect 8568 5326 8602 5328
rect -96 5298 -54 5300
rect 1238 5298 1272 5300
rect 4886 5298 4928 5300
rect 6220 5298 6254 5300
rect 7908 4712 7982 4740
rect 7908 4700 7926 4712
rect 7960 4700 7982 4712
rect 7908 4496 7982 4516
rect 7908 4462 7926 4496
rect 7960 4462 7982 4496
rect 7908 4452 7982 4462
rect 7926 4432 7960 4452
rect 7714 4278 7778 4296
rect 7962 4278 8002 4296
rect 7694 4244 7724 4278
rect 7758 4244 7778 4278
rect 7974 4244 8002 4278
rect 7714 4222 7778 4244
rect 7962 4222 8002 4244
rect 8150 3154 8210 3190
rect 9074 3154 9160 3190
rect 8154 3054 8164 3088
rect 8198 3054 8214 3088
rect 9078 3054 9100 3088
rect 9134 3054 9164 3088
rect 8154 3052 8214 3054
rect 9078 3052 9164 3054
rect 8156 2960 8166 2994
rect 8200 2960 8216 2994
rect 9080 2960 9102 2994
rect 9136 2960 9166 2994
rect 8156 2958 8216 2960
rect 9080 2958 9166 2960
rect 8156 2848 8166 2882
rect 8200 2848 8216 2882
rect 9080 2848 9102 2882
rect 9136 2848 9166 2882
rect 8156 2846 8216 2848
rect 9080 2846 9166 2848
rect 7708 2732 7768 2734
rect 9136 2732 9182 2734
rect -440 2714 -380 2716
rect 988 2714 1034 2716
rect -3072 2704 -3012 2706
rect -1644 2704 -1598 2706
rect -4962 2652 -4902 2692
rect -3534 2652 -3488 2692
rect -3072 2670 -3040 2704
rect -1638 2670 -1598 2704
rect -440 2680 -408 2714
rect 994 2680 1034 2714
rect -440 2676 -380 2680
rect 988 2676 1034 2680
rect 2298 2704 2358 2706
rect 3726 2704 3772 2706
rect -3072 2666 -3012 2670
rect -1644 2666 -1598 2670
rect 2298 2670 2330 2704
rect 3732 2670 3772 2704
rect 7708 2698 7740 2732
rect 9142 2698 9182 2732
rect 7708 2694 7768 2698
rect 9136 2694 9182 2698
rect 2298 2666 2358 2670
rect 3726 2666 3772 2670
rect 4998 2676 5058 2678
rect 6426 2676 6472 2678
rect 4998 2642 5030 2676
rect 6432 2642 6472 2676
rect 4998 2638 5058 2642
rect 6426 2638 6472 2642
rect 7706 2632 7766 2638
rect 9134 2632 9180 2638
rect -442 2614 -382 2620
rect 986 2614 1032 2620
rect -3074 2604 -3014 2610
rect -1646 2604 -1600 2610
rect -4964 2556 -4904 2596
rect -3536 2556 -3490 2596
rect -3074 2570 -3040 2604
rect -1638 2570 -1600 2604
rect -442 2580 -408 2614
rect 994 2580 1032 2614
rect 2296 2604 2356 2610
rect 3724 2604 3770 2610
rect 2296 2570 2330 2604
rect 3732 2570 3770 2604
rect 7706 2598 7740 2632
rect 9142 2598 9180 2632
rect 4996 2576 5056 2582
rect 6424 2576 6470 2582
rect 4996 2542 5030 2576
rect 6432 2542 6470 2576
<< viali >>
rect -2710 5410 -2682 5444
rect -2682 5410 -2676 5444
rect -2638 5410 -2604 5444
rect -2566 5410 -2532 5444
rect -2494 5410 -2460 5444
rect -2422 5410 -2388 5444
rect -2350 5410 -2316 5444
rect -2278 5410 -2244 5444
rect -2206 5410 -2172 5444
rect -2134 5410 -2100 5444
rect -2062 5410 -2028 5444
rect -1990 5410 -1956 5444
rect -1918 5410 -1884 5444
rect -1846 5410 -1812 5444
rect -1774 5410 -1740 5444
rect -1702 5410 -1668 5444
rect -1630 5410 -1596 5444
rect -1558 5410 -1524 5444
rect -1486 5410 -1452 5444
rect -1414 5410 -1390 5444
rect -1390 5410 -1380 5444
rect -1342 5410 -1308 5444
rect -78 5400 -50 5434
rect -50 5400 -44 5434
rect -6 5400 28 5434
rect 66 5400 100 5434
rect 138 5400 172 5434
rect 210 5400 244 5434
rect 282 5400 316 5434
rect 354 5400 388 5434
rect 426 5400 460 5434
rect 498 5400 532 5434
rect 570 5400 604 5434
rect 642 5400 676 5434
rect 714 5400 748 5434
rect 786 5400 820 5434
rect 858 5400 892 5434
rect 930 5400 964 5434
rect 1002 5400 1036 5434
rect 1074 5400 1108 5434
rect 1146 5400 1180 5434
rect 1218 5400 1242 5434
rect 1242 5400 1252 5434
rect 1290 5400 1324 5434
rect 2280 5428 2308 5462
rect 2308 5428 2314 5462
rect 2352 5428 2386 5462
rect 2424 5428 2458 5462
rect 2496 5428 2530 5462
rect 2568 5428 2602 5462
rect 2640 5428 2674 5462
rect 2712 5428 2746 5462
rect 2784 5428 2818 5462
rect 2856 5428 2890 5462
rect 2928 5428 2962 5462
rect 3000 5428 3034 5462
rect 3072 5428 3106 5462
rect 3144 5428 3178 5462
rect 3216 5428 3250 5462
rect 3288 5428 3322 5462
rect 3360 5428 3394 5462
rect 3432 5428 3466 5462
rect 3504 5428 3538 5462
rect 3576 5428 3600 5462
rect 3600 5428 3610 5462
rect 3648 5428 3682 5462
rect 4904 5400 4932 5434
rect 4932 5400 4938 5434
rect 4976 5400 5010 5434
rect 5048 5400 5082 5434
rect 5120 5400 5154 5434
rect 5192 5400 5226 5434
rect 5264 5400 5298 5434
rect 5336 5400 5370 5434
rect 5408 5400 5442 5434
rect 5480 5400 5514 5434
rect 5552 5400 5586 5434
rect 5624 5400 5658 5434
rect 5696 5400 5730 5434
rect 5768 5400 5802 5434
rect 5840 5400 5874 5434
rect 5912 5400 5946 5434
rect 5984 5400 6018 5434
rect 6056 5400 6090 5434
rect 6128 5400 6162 5434
rect 6200 5400 6224 5434
rect 6224 5400 6234 5434
rect 6272 5400 6306 5434
rect 7252 5428 7280 5462
rect 7280 5428 7286 5462
rect 7324 5428 7358 5462
rect 7396 5428 7430 5462
rect 7468 5428 7502 5462
rect 7540 5428 7574 5462
rect 7612 5428 7646 5462
rect 7684 5428 7718 5462
rect 7756 5428 7790 5462
rect 7828 5428 7862 5462
rect 7900 5428 7934 5462
rect 7972 5428 8006 5462
rect 8044 5428 8078 5462
rect 8116 5428 8150 5462
rect 8188 5428 8222 5462
rect 8260 5428 8294 5462
rect 8332 5428 8366 5462
rect 8404 5428 8438 5462
rect 8476 5428 8510 5462
rect 8548 5428 8572 5462
rect 8572 5428 8582 5462
rect 8620 5428 8654 5462
rect -2718 5310 -2686 5344
rect -2686 5310 -2684 5344
rect -2646 5310 -2612 5344
rect -2574 5310 -2540 5344
rect -2502 5310 -2468 5344
rect -2430 5310 -2396 5344
rect -2358 5310 -2324 5344
rect -2286 5310 -2252 5344
rect -2214 5310 -2180 5344
rect -2142 5310 -2108 5344
rect -2070 5310 -2036 5344
rect -1998 5310 -1964 5344
rect -1926 5310 -1892 5344
rect -1854 5310 -1820 5344
rect -1782 5310 -1748 5344
rect -1710 5310 -1676 5344
rect -1638 5310 -1604 5344
rect -1566 5310 -1532 5344
rect -1494 5310 -1460 5344
rect -1422 5310 -1394 5344
rect -1394 5310 -1388 5344
rect -1350 5310 -1316 5344
rect -86 5300 -54 5334
rect -54 5300 -52 5334
rect -14 5300 20 5334
rect 58 5300 92 5334
rect 130 5300 164 5334
rect 202 5300 236 5334
rect 274 5300 308 5334
rect 346 5300 380 5334
rect 418 5300 452 5334
rect 490 5300 524 5334
rect 562 5300 596 5334
rect 634 5300 668 5334
rect 706 5300 740 5334
rect 778 5300 812 5334
rect 850 5300 884 5334
rect 922 5300 956 5334
rect 994 5300 1028 5334
rect 1066 5300 1100 5334
rect 1138 5300 1172 5334
rect 1210 5300 1238 5334
rect 1238 5300 1244 5334
rect 1282 5300 1316 5334
rect 2272 5328 2304 5362
rect 2304 5328 2306 5362
rect 2344 5328 2378 5362
rect 2416 5328 2450 5362
rect 2488 5328 2522 5362
rect 2560 5328 2594 5362
rect 2632 5328 2666 5362
rect 2704 5328 2738 5362
rect 2776 5328 2810 5362
rect 2848 5328 2882 5362
rect 2920 5328 2954 5362
rect 2992 5328 3026 5362
rect 3064 5328 3098 5362
rect 3136 5328 3170 5362
rect 3208 5328 3242 5362
rect 3280 5328 3314 5362
rect 3352 5328 3386 5362
rect 3424 5328 3458 5362
rect 3496 5328 3530 5362
rect 3568 5328 3596 5362
rect 3596 5328 3602 5362
rect 3640 5328 3674 5362
rect 4896 5300 4928 5334
rect 4928 5300 4930 5334
rect 4968 5300 5002 5334
rect 5040 5300 5074 5334
rect 5112 5300 5146 5334
rect 5184 5300 5218 5334
rect 5256 5300 5290 5334
rect 5328 5300 5362 5334
rect 5400 5300 5434 5334
rect 5472 5300 5506 5334
rect 5544 5300 5578 5334
rect 5616 5300 5650 5334
rect 5688 5300 5722 5334
rect 5760 5300 5794 5334
rect 5832 5300 5866 5334
rect 5904 5300 5938 5334
rect 5976 5300 6010 5334
rect 6048 5300 6082 5334
rect 6120 5300 6154 5334
rect 6192 5300 6220 5334
rect 6220 5300 6226 5334
rect 6264 5300 6298 5334
rect 7244 5328 7276 5362
rect 7276 5328 7278 5362
rect 7316 5328 7350 5362
rect 7388 5328 7422 5362
rect 7460 5328 7494 5362
rect 7532 5328 7566 5362
rect 7604 5328 7638 5362
rect 7676 5328 7710 5362
rect 7748 5328 7782 5362
rect 7820 5328 7854 5362
rect 7892 5328 7926 5362
rect 7964 5328 7998 5362
rect 8036 5328 8070 5362
rect 8108 5328 8142 5362
rect 8180 5328 8214 5362
rect 8252 5328 8286 5362
rect 8324 5328 8358 5362
rect 8396 5328 8430 5362
rect 8468 5328 8502 5362
rect 8540 5328 8568 5362
rect 8568 5328 8574 5362
rect 8612 5328 8646 5362
rect 7926 4700 7960 4712
rect 7926 4678 7960 4700
rect 7926 4606 7960 4640
rect 7926 4534 7960 4568
rect 7926 4462 7960 4496
rect 7724 4244 7758 4278
rect 7796 4244 7830 4278
rect 7868 4244 7902 4278
rect 7940 4244 7962 4278
rect 7962 4244 7974 4278
rect -3792 4050 -3742 4108
rect -4398 3878 -4348 3936
rect 8538 3876 8588 3934
rect 8164 3054 8198 3088
rect 8236 3054 8270 3088
rect 8308 3054 8342 3088
rect 8380 3054 8414 3088
rect 8452 3054 8486 3088
rect 8524 3054 8558 3088
rect 8596 3054 8630 3088
rect 8668 3054 8702 3088
rect 8740 3054 8774 3088
rect 8812 3054 8846 3088
rect 8884 3054 8918 3088
rect 8956 3054 8990 3088
rect 9028 3054 9062 3088
rect 9100 3054 9134 3088
rect 8166 2960 8200 2994
rect 8238 2960 8272 2994
rect 8310 2960 8344 2994
rect 8382 2960 8416 2994
rect 8454 2960 8488 2994
rect 8526 2960 8560 2994
rect 8598 2960 8632 2994
rect 8670 2960 8704 2994
rect 8742 2960 8776 2994
rect 8814 2960 8848 2994
rect 8886 2960 8920 2994
rect 8958 2960 8992 2994
rect 9030 2960 9064 2994
rect 9102 2960 9136 2994
rect 8166 2848 8200 2882
rect 8238 2848 8272 2882
rect 8310 2848 8344 2882
rect 8382 2848 8416 2882
rect 8454 2848 8488 2882
rect 8526 2848 8560 2882
rect 8598 2848 8632 2882
rect 8670 2848 8704 2882
rect 8742 2848 8776 2882
rect 8814 2848 8848 2882
rect 8886 2848 8920 2882
rect 8958 2848 8992 2882
rect 9030 2848 9064 2882
rect 9102 2848 9136 2882
rect -3040 2670 -3012 2704
rect -3012 2670 -3006 2704
rect -2968 2670 -2934 2704
rect -2896 2670 -2862 2704
rect -2824 2670 -2790 2704
rect -2752 2670 -2718 2704
rect -2680 2670 -2646 2704
rect -2608 2670 -2574 2704
rect -2536 2670 -2502 2704
rect -2464 2670 -2430 2704
rect -2392 2670 -2358 2704
rect -2320 2670 -2286 2704
rect -2248 2670 -2214 2704
rect -2176 2670 -2142 2704
rect -2104 2670 -2070 2704
rect -2032 2670 -1998 2704
rect -1960 2670 -1926 2704
rect -1888 2670 -1854 2704
rect -1816 2670 -1782 2704
rect -1744 2670 -1710 2704
rect -1672 2670 -1644 2704
rect -1644 2670 -1638 2704
rect -408 2680 -380 2714
rect -380 2680 -374 2714
rect -336 2680 -302 2714
rect -264 2680 -230 2714
rect -192 2680 -158 2714
rect -120 2680 -86 2714
rect -48 2680 -14 2714
rect 24 2680 58 2714
rect 96 2680 130 2714
rect 168 2680 202 2714
rect 240 2680 274 2714
rect 312 2680 346 2714
rect 384 2680 418 2714
rect 456 2680 490 2714
rect 528 2680 562 2714
rect 600 2680 634 2714
rect 672 2680 706 2714
rect 744 2680 778 2714
rect 816 2680 850 2714
rect 888 2680 922 2714
rect 960 2680 988 2714
rect 988 2680 994 2714
rect 2330 2670 2358 2704
rect 2358 2670 2364 2704
rect 2402 2670 2436 2704
rect 2474 2670 2508 2704
rect 2546 2670 2580 2704
rect 2618 2670 2652 2704
rect 2690 2670 2724 2704
rect 2762 2670 2796 2704
rect 2834 2670 2868 2704
rect 2906 2670 2940 2704
rect 2978 2670 3012 2704
rect 3050 2670 3084 2704
rect 3122 2670 3156 2704
rect 3194 2670 3228 2704
rect 3266 2670 3300 2704
rect 3338 2670 3372 2704
rect 3410 2670 3444 2704
rect 3482 2670 3516 2704
rect 3554 2670 3588 2704
rect 3626 2670 3660 2704
rect 3698 2670 3726 2704
rect 3726 2670 3732 2704
rect 7740 2698 7768 2732
rect 7768 2698 7774 2732
rect 7812 2698 7846 2732
rect 7884 2698 7918 2732
rect 7956 2698 7990 2732
rect 8028 2698 8062 2732
rect 8100 2698 8134 2732
rect 8172 2698 8206 2732
rect 8244 2698 8278 2732
rect 8316 2698 8350 2732
rect 8388 2698 8422 2732
rect 8460 2698 8494 2732
rect 8532 2698 8566 2732
rect 8604 2698 8638 2732
rect 8676 2698 8710 2732
rect 8748 2698 8782 2732
rect 8820 2698 8854 2732
rect 8892 2698 8926 2732
rect 8964 2698 8998 2732
rect 9036 2698 9070 2732
rect 9108 2698 9136 2732
rect 9136 2698 9142 2732
rect 5030 2642 5058 2676
rect 5058 2642 5064 2676
rect 5102 2642 5136 2676
rect 5174 2642 5208 2676
rect 5246 2642 5280 2676
rect 5318 2642 5352 2676
rect 5390 2642 5424 2676
rect 5462 2642 5496 2676
rect 5534 2642 5568 2676
rect 5606 2642 5640 2676
rect 5678 2642 5712 2676
rect 5750 2642 5784 2676
rect 5822 2642 5856 2676
rect 5894 2642 5928 2676
rect 5966 2642 6000 2676
rect 6038 2642 6072 2676
rect 6110 2642 6144 2676
rect 6182 2642 6216 2676
rect 6254 2642 6288 2676
rect 6326 2642 6360 2676
rect 6398 2642 6426 2676
rect 6426 2642 6432 2676
rect -3040 2570 -3014 2604
rect -3014 2570 -3006 2604
rect -2968 2570 -2934 2604
rect -2896 2570 -2862 2604
rect -2824 2570 -2790 2604
rect -2752 2570 -2718 2604
rect -2680 2570 -2646 2604
rect -2608 2570 -2574 2604
rect -2536 2570 -2502 2604
rect -2464 2570 -2430 2604
rect -2392 2570 -2358 2604
rect -2320 2570 -2286 2604
rect -2248 2570 -2214 2604
rect -2176 2570 -2142 2604
rect -2104 2570 -2070 2604
rect -2032 2570 -1998 2604
rect -1960 2570 -1926 2604
rect -1888 2570 -1854 2604
rect -1816 2570 -1782 2604
rect -1744 2570 -1710 2604
rect -1672 2570 -1646 2604
rect -1646 2570 -1638 2604
rect -408 2580 -382 2614
rect -382 2580 -374 2614
rect -336 2580 -302 2614
rect -264 2580 -230 2614
rect -192 2580 -158 2614
rect -120 2580 -86 2614
rect -48 2580 -14 2614
rect 24 2580 58 2614
rect 96 2580 130 2614
rect 168 2580 202 2614
rect 240 2580 274 2614
rect 312 2580 346 2614
rect 384 2580 418 2614
rect 456 2580 490 2614
rect 528 2580 562 2614
rect 600 2580 634 2614
rect 672 2580 706 2614
rect 744 2580 778 2614
rect 816 2580 850 2614
rect 888 2580 922 2614
rect 960 2580 986 2614
rect 986 2580 994 2614
rect 2330 2570 2356 2604
rect 2356 2570 2364 2604
rect 2402 2570 2436 2604
rect 2474 2570 2508 2604
rect 2546 2570 2580 2604
rect 2618 2570 2652 2604
rect 2690 2570 2724 2604
rect 2762 2570 2796 2604
rect 2834 2570 2868 2604
rect 2906 2570 2940 2604
rect 2978 2570 3012 2604
rect 3050 2570 3084 2604
rect 3122 2570 3156 2604
rect 3194 2570 3228 2604
rect 3266 2570 3300 2604
rect 3338 2570 3372 2604
rect 3410 2570 3444 2604
rect 3482 2570 3516 2604
rect 3554 2570 3588 2604
rect 3626 2570 3660 2604
rect 3698 2570 3724 2604
rect 3724 2570 3732 2604
rect 7740 2598 7766 2632
rect 7766 2598 7774 2632
rect 7812 2598 7846 2632
rect 7884 2598 7918 2632
rect 7956 2598 7990 2632
rect 8028 2598 8062 2632
rect 8100 2598 8134 2632
rect 8172 2598 8206 2632
rect 8244 2598 8278 2632
rect 8316 2598 8350 2632
rect 8388 2598 8422 2632
rect 8460 2598 8494 2632
rect 8532 2598 8566 2632
rect 8604 2598 8638 2632
rect 8676 2598 8710 2632
rect 8748 2598 8782 2632
rect 8820 2598 8854 2632
rect 8892 2598 8926 2632
rect 8964 2598 8998 2632
rect 9036 2598 9070 2632
rect 9108 2598 9134 2632
rect 9134 2598 9142 2632
rect 5030 2542 5056 2576
rect 5056 2542 5064 2576
rect 5102 2542 5136 2576
rect 5174 2542 5208 2576
rect 5246 2542 5280 2576
rect 5318 2542 5352 2576
rect 5390 2542 5424 2576
rect 5462 2542 5496 2576
rect 5534 2542 5568 2576
rect 5606 2542 5640 2576
rect 5678 2542 5712 2576
rect 5750 2542 5784 2576
rect 5822 2542 5856 2576
rect 5894 2542 5928 2576
rect 5966 2542 6000 2576
rect 6038 2542 6072 2576
rect 6110 2542 6144 2576
rect 6182 2542 6216 2576
rect 6254 2542 6288 2576
rect 6326 2542 6360 2576
rect 6398 2542 6424 2576
rect 6424 2542 6432 2576
<< metal1 >>
rect -5122 5462 9233 5516
rect -5122 5444 2280 5462
rect -5122 5410 -2710 5444
rect -2676 5410 -2638 5444
rect -2604 5410 -2566 5444
rect -2532 5410 -2494 5444
rect -2460 5410 -2422 5444
rect -2388 5410 -2350 5444
rect -2316 5410 -2278 5444
rect -2244 5410 -2206 5444
rect -2172 5410 -2134 5444
rect -2100 5410 -2062 5444
rect -2028 5410 -1990 5444
rect -1956 5410 -1918 5444
rect -1884 5410 -1846 5444
rect -1812 5410 -1774 5444
rect -1740 5410 -1702 5444
rect -1668 5410 -1630 5444
rect -1596 5410 -1558 5444
rect -1524 5410 -1486 5444
rect -1452 5410 -1414 5444
rect -1380 5410 -1342 5444
rect -1308 5434 2280 5444
rect -1308 5410 -78 5434
rect -5122 5400 -78 5410
rect -44 5400 -6 5434
rect 28 5400 66 5434
rect 100 5400 138 5434
rect 172 5400 210 5434
rect 244 5400 282 5434
rect 316 5400 354 5434
rect 388 5400 426 5434
rect 460 5400 498 5434
rect 532 5400 570 5434
rect 604 5400 642 5434
rect 676 5400 714 5434
rect 748 5400 786 5434
rect 820 5400 858 5434
rect 892 5400 930 5434
rect 964 5400 1002 5434
rect 1036 5400 1074 5434
rect 1108 5400 1146 5434
rect 1180 5400 1218 5434
rect 1252 5400 1290 5434
rect 1324 5428 2280 5434
rect 2314 5428 2352 5462
rect 2386 5428 2424 5462
rect 2458 5428 2496 5462
rect 2530 5428 2568 5462
rect 2602 5428 2640 5462
rect 2674 5428 2712 5462
rect 2746 5428 2784 5462
rect 2818 5428 2856 5462
rect 2890 5428 2928 5462
rect 2962 5428 3000 5462
rect 3034 5428 3072 5462
rect 3106 5428 3144 5462
rect 3178 5428 3216 5462
rect 3250 5428 3288 5462
rect 3322 5428 3360 5462
rect 3394 5428 3432 5462
rect 3466 5428 3504 5462
rect 3538 5428 3576 5462
rect 3610 5428 3648 5462
rect 3682 5434 7252 5462
rect 3682 5428 4904 5434
rect 1324 5400 4904 5428
rect 4938 5400 4976 5434
rect 5010 5400 5048 5434
rect 5082 5400 5120 5434
rect 5154 5400 5192 5434
rect 5226 5400 5264 5434
rect 5298 5400 5336 5434
rect 5370 5400 5408 5434
rect 5442 5400 5480 5434
rect 5514 5400 5552 5434
rect 5586 5400 5624 5434
rect 5658 5400 5696 5434
rect 5730 5400 5768 5434
rect 5802 5400 5840 5434
rect 5874 5400 5912 5434
rect 5946 5400 5984 5434
rect 6018 5400 6056 5434
rect 6090 5400 6128 5434
rect 6162 5400 6200 5434
rect 6234 5400 6272 5434
rect 6306 5428 7252 5434
rect 7286 5428 7324 5462
rect 7358 5428 7396 5462
rect 7430 5428 7468 5462
rect 7502 5428 7540 5462
rect 7574 5428 7612 5462
rect 7646 5428 7684 5462
rect 7718 5428 7756 5462
rect 7790 5428 7828 5462
rect 7862 5428 7900 5462
rect 7934 5428 7972 5462
rect 8006 5428 8044 5462
rect 8078 5428 8116 5462
rect 8150 5428 8188 5462
rect 8222 5428 8260 5462
rect 8294 5428 8332 5462
rect 8366 5428 8404 5462
rect 8438 5428 8476 5462
rect 8510 5428 8548 5462
rect 8582 5428 8620 5462
rect 8654 5428 9233 5462
rect 6306 5400 9233 5428
rect -5122 5362 9233 5400
rect -5122 5344 2272 5362
rect -5122 5310 -2718 5344
rect -2684 5310 -2646 5344
rect -2612 5310 -2574 5344
rect -2540 5310 -2502 5344
rect -2468 5310 -2430 5344
rect -2396 5310 -2358 5344
rect -2324 5310 -2286 5344
rect -2252 5310 -2214 5344
rect -2180 5310 -2142 5344
rect -2108 5310 -2070 5344
rect -2036 5310 -1998 5344
rect -1964 5310 -1926 5344
rect -1892 5310 -1854 5344
rect -1820 5310 -1782 5344
rect -1748 5310 -1710 5344
rect -1676 5310 -1638 5344
rect -1604 5310 -1566 5344
rect -1532 5310 -1494 5344
rect -1460 5310 -1422 5344
rect -1388 5310 -1350 5344
rect -1316 5334 2272 5344
rect -1316 5310 -86 5334
rect -5122 5300 -86 5310
rect -52 5300 -14 5334
rect 20 5300 58 5334
rect 92 5300 130 5334
rect 164 5300 202 5334
rect 236 5300 274 5334
rect 308 5300 346 5334
rect 380 5300 418 5334
rect 452 5300 490 5334
rect 524 5300 562 5334
rect 596 5300 634 5334
rect 668 5300 706 5334
rect 740 5300 778 5334
rect 812 5300 850 5334
rect 884 5300 922 5334
rect 956 5300 994 5334
rect 1028 5300 1066 5334
rect 1100 5300 1138 5334
rect 1172 5300 1210 5334
rect 1244 5300 1282 5334
rect 1316 5328 2272 5334
rect 2306 5328 2344 5362
rect 2378 5328 2416 5362
rect 2450 5328 2488 5362
rect 2522 5328 2560 5362
rect 2594 5328 2632 5362
rect 2666 5328 2704 5362
rect 2738 5328 2776 5362
rect 2810 5328 2848 5362
rect 2882 5328 2920 5362
rect 2954 5328 2992 5362
rect 3026 5328 3064 5362
rect 3098 5328 3136 5362
rect 3170 5328 3208 5362
rect 3242 5328 3280 5362
rect 3314 5328 3352 5362
rect 3386 5328 3424 5362
rect 3458 5328 3496 5362
rect 3530 5328 3568 5362
rect 3602 5328 3640 5362
rect 3674 5334 7244 5362
rect 3674 5328 4896 5334
rect 1316 5300 4896 5328
rect 4930 5300 4968 5334
rect 5002 5300 5040 5334
rect 5074 5300 5112 5334
rect 5146 5300 5184 5334
rect 5218 5300 5256 5334
rect 5290 5300 5328 5334
rect 5362 5300 5400 5334
rect 5434 5300 5472 5334
rect 5506 5300 5544 5334
rect 5578 5300 5616 5334
rect 5650 5300 5688 5334
rect 5722 5300 5760 5334
rect 5794 5300 5832 5334
rect 5866 5300 5904 5334
rect 5938 5300 5976 5334
rect 6010 5300 6048 5334
rect 6082 5300 6120 5334
rect 6154 5300 6192 5334
rect 6226 5300 6264 5334
rect 6298 5328 7244 5334
rect 7278 5328 7316 5362
rect 7350 5328 7388 5362
rect 7422 5328 7460 5362
rect 7494 5328 7532 5362
rect 7566 5328 7604 5362
rect 7638 5328 7676 5362
rect 7710 5328 7748 5362
rect 7782 5328 7820 5362
rect 7854 5328 7892 5362
rect 7926 5328 7964 5362
rect 7998 5328 8036 5362
rect 8070 5328 8108 5362
rect 8142 5328 8180 5362
rect 8214 5328 8252 5362
rect 8286 5328 8324 5362
rect 8358 5328 8396 5362
rect 8430 5328 8468 5362
rect 8502 5328 8540 5362
rect 8574 5328 8612 5362
rect 8646 5328 9233 5362
rect 6298 5300 9233 5328
rect -5122 5198 9233 5300
rect -4874 5051 -4832 5198
rect -4804 5082 -4794 5142
rect -4734 5082 -4724 5142
rect -4874 4888 -4790 5051
rect -3768 5046 -3726 5198
rect -3698 5088 -3688 5148
rect -3628 5088 -3618 5148
rect -4726 5040 -4470 5046
rect -4736 5032 -4470 5040
rect -4874 4886 -4832 4888
rect -4740 4882 -4730 5032
rect -4674 4882 -4470 5032
rect -4896 3112 -4822 3114
rect -4898 2932 -4822 3112
rect -4736 3109 -4470 4882
rect -3768 4849 -3698 5046
rect -3636 4352 -3499 5046
rect 7850 4712 8202 4866
rect 7850 4678 7926 4712
rect 7960 4678 8202 4712
rect 7850 4640 8202 4678
rect 7850 4606 7926 4640
rect 7960 4606 8202 4640
rect 7850 4568 8202 4606
rect 8741 4706 9233 5198
rect 7850 4534 7926 4568
rect 7960 4534 8202 4568
rect 7850 4496 8202 4534
rect 7850 4462 7926 4496
rect 7960 4462 8202 4496
rect 7850 4352 8202 4462
rect -4314 4278 8202 4352
rect -4314 4244 7724 4278
rect 7758 4244 7796 4278
rect 7830 4244 7868 4278
rect 7902 4244 7940 4278
rect 7974 4244 8202 4278
rect -4314 4172 8202 4244
rect -3798 4108 -3736 4120
rect -3798 4050 -3792 4108
rect -3742 4050 -3736 4108
rect -3798 4038 -3736 4050
rect -4404 3936 -4342 3948
rect -4404 3878 -4398 3936
rect -4348 3878 -4342 3936
rect -4404 3866 -4342 3878
rect 8258 3922 8292 4592
rect 8741 4451 9231 4706
rect 8960 4160 8994 4451
rect 8532 3934 8594 3946
rect 8532 3922 8538 3934
rect 8258 3886 8538 3922
rect 8168 3624 8202 3684
rect -4767 2937 -4470 3109
rect -3770 2956 -3696 3138
rect -4736 2935 -4470 2937
rect -4898 2804 -4862 2932
rect -4834 2848 -4824 2902
rect -4764 2848 -4754 2902
rect -3768 2804 -3732 2956
rect -3640 2950 -3608 3532
rect 7804 3520 8202 3624
rect 8168 3444 8202 3520
rect 8258 3474 8292 3886
rect 8532 3876 8538 3886
rect 8588 3922 8594 3934
rect 8588 3920 8689 3922
rect 9050 3920 9082 4350
rect 8588 3886 8693 3920
rect 9050 3886 9347 3920
rect 8588 3876 8594 3886
rect 8532 3864 8594 3876
rect 8343 3351 8400 3419
rect 8960 3417 8996 3620
rect 9050 3526 9082 3886
rect 8092 3220 8400 3351
rect 8602 3220 9243 3417
rect 8093 3088 9245 3220
rect 8093 3054 8164 3088
rect 8198 3054 8236 3088
rect 8270 3054 8308 3088
rect 8342 3054 8380 3088
rect 8414 3054 8452 3088
rect 8486 3054 8524 3088
rect 8558 3054 8596 3088
rect 8630 3054 8668 3088
rect 8702 3054 8740 3088
rect 8774 3054 8812 3088
rect 8846 3054 8884 3088
rect 8918 3054 8956 3088
rect 8990 3054 9028 3088
rect 9062 3054 9100 3088
rect 9134 3054 9245 3088
rect 8093 2994 9245 3054
rect 8093 2960 8166 2994
rect 8200 2960 8238 2994
rect 8272 2960 8310 2994
rect 8344 2960 8382 2994
rect 8416 2960 8454 2994
rect 8488 2960 8526 2994
rect 8560 2960 8598 2994
rect 8632 2960 8670 2994
rect 8704 2960 8742 2994
rect 8776 2960 8814 2994
rect 8848 2960 8886 2994
rect 8920 2960 8958 2994
rect 8992 2960 9030 2994
rect 9064 2960 9102 2994
rect 9136 2960 9245 2994
rect -3702 2844 -3692 2898
rect -3632 2844 -3622 2898
rect 8093 2882 9245 2960
rect 8093 2848 8166 2882
rect 8200 2848 8238 2882
rect 8272 2848 8310 2882
rect 8344 2848 8382 2882
rect 8416 2848 8454 2882
rect 8488 2848 8526 2882
rect 8560 2848 8598 2882
rect 8632 2848 8670 2882
rect 8704 2848 8742 2882
rect 8776 2848 8814 2882
rect 8848 2848 8886 2882
rect 8920 2848 8958 2882
rect 8992 2848 9030 2882
rect 9064 2848 9102 2882
rect 9136 2848 9245 2882
rect 8093 2804 9245 2848
rect -5118 2732 9245 2804
rect -5118 2714 7740 2732
rect -5118 2704 -408 2714
rect -5118 2670 -3040 2704
rect -3006 2670 -2968 2704
rect -2934 2670 -2896 2704
rect -2862 2670 -2824 2704
rect -2790 2670 -2752 2704
rect -2718 2670 -2680 2704
rect -2646 2670 -2608 2704
rect -2574 2670 -2536 2704
rect -2502 2670 -2464 2704
rect -2430 2670 -2392 2704
rect -2358 2670 -2320 2704
rect -2286 2670 -2248 2704
rect -2214 2670 -2176 2704
rect -2142 2670 -2104 2704
rect -2070 2670 -2032 2704
rect -1998 2670 -1960 2704
rect -1926 2670 -1888 2704
rect -1854 2670 -1816 2704
rect -1782 2670 -1744 2704
rect -1710 2670 -1672 2704
rect -1638 2680 -408 2704
rect -374 2680 -336 2714
rect -302 2680 -264 2714
rect -230 2680 -192 2714
rect -158 2680 -120 2714
rect -86 2680 -48 2714
rect -14 2680 24 2714
rect 58 2680 96 2714
rect 130 2680 168 2714
rect 202 2680 240 2714
rect 274 2680 312 2714
rect 346 2680 384 2714
rect 418 2680 456 2714
rect 490 2680 528 2714
rect 562 2680 600 2714
rect 634 2680 672 2714
rect 706 2680 744 2714
rect 778 2680 816 2714
rect 850 2680 888 2714
rect 922 2680 960 2714
rect 994 2704 7740 2714
rect 994 2680 2330 2704
rect -1638 2670 2330 2680
rect 2364 2670 2402 2704
rect 2436 2670 2474 2704
rect 2508 2670 2546 2704
rect 2580 2670 2618 2704
rect 2652 2670 2690 2704
rect 2724 2670 2762 2704
rect 2796 2670 2834 2704
rect 2868 2670 2906 2704
rect 2940 2670 2978 2704
rect 3012 2670 3050 2704
rect 3084 2670 3122 2704
rect 3156 2670 3194 2704
rect 3228 2670 3266 2704
rect 3300 2670 3338 2704
rect 3372 2670 3410 2704
rect 3444 2670 3482 2704
rect 3516 2670 3554 2704
rect 3588 2670 3626 2704
rect 3660 2670 3698 2704
rect 3732 2698 7740 2704
rect 7774 2698 7812 2732
rect 7846 2698 7884 2732
rect 7918 2698 7956 2732
rect 7990 2698 8028 2732
rect 8062 2698 8100 2732
rect 8134 2698 8172 2732
rect 8206 2698 8244 2732
rect 8278 2698 8316 2732
rect 8350 2698 8388 2732
rect 8422 2698 8460 2732
rect 8494 2698 8532 2732
rect 8566 2698 8604 2732
rect 8638 2698 8676 2732
rect 8710 2698 8748 2732
rect 8782 2698 8820 2732
rect 8854 2698 8892 2732
rect 8926 2698 8964 2732
rect 8998 2698 9036 2732
rect 9070 2698 9108 2732
rect 9142 2698 9245 2732
rect 3732 2676 9245 2698
rect 3732 2670 5030 2676
rect -5118 2642 5030 2670
rect 5064 2642 5102 2676
rect 5136 2642 5174 2676
rect 5208 2642 5246 2676
rect 5280 2642 5318 2676
rect 5352 2642 5390 2676
rect 5424 2642 5462 2676
rect 5496 2642 5534 2676
rect 5568 2642 5606 2676
rect 5640 2642 5678 2676
rect 5712 2642 5750 2676
rect 5784 2642 5822 2676
rect 5856 2642 5894 2676
rect 5928 2642 5966 2676
rect 6000 2642 6038 2676
rect 6072 2642 6110 2676
rect 6144 2642 6182 2676
rect 6216 2642 6254 2676
rect 6288 2642 6326 2676
rect 6360 2642 6398 2676
rect 6432 2642 9245 2676
rect -5118 2632 9245 2642
rect -5118 2624 7740 2632
rect -5114 2614 7740 2624
rect -5114 2604 -408 2614
rect -5114 2570 -3040 2604
rect -3006 2570 -2968 2604
rect -2934 2570 -2896 2604
rect -2862 2570 -2824 2604
rect -2790 2570 -2752 2604
rect -2718 2570 -2680 2604
rect -2646 2570 -2608 2604
rect -2574 2570 -2536 2604
rect -2502 2570 -2464 2604
rect -2430 2570 -2392 2604
rect -2358 2570 -2320 2604
rect -2286 2570 -2248 2604
rect -2214 2570 -2176 2604
rect -2142 2570 -2104 2604
rect -2070 2570 -2032 2604
rect -1998 2570 -1960 2604
rect -1926 2570 -1888 2604
rect -1854 2570 -1816 2604
rect -1782 2570 -1744 2604
rect -1710 2570 -1672 2604
rect -1638 2580 -408 2604
rect -374 2580 -336 2614
rect -302 2580 -264 2614
rect -230 2580 -192 2614
rect -158 2580 -120 2614
rect -86 2580 -48 2614
rect -14 2580 24 2614
rect 58 2580 96 2614
rect 130 2580 168 2614
rect 202 2580 240 2614
rect 274 2580 312 2614
rect 346 2580 384 2614
rect 418 2580 456 2614
rect 490 2580 528 2614
rect 562 2580 600 2614
rect 634 2580 672 2614
rect 706 2580 744 2614
rect 778 2580 816 2614
rect 850 2580 888 2614
rect 922 2580 960 2614
rect 994 2604 7740 2614
rect 994 2580 2330 2604
rect -1638 2570 2330 2580
rect 2364 2570 2402 2604
rect 2436 2570 2474 2604
rect 2508 2570 2546 2604
rect 2580 2570 2618 2604
rect 2652 2570 2690 2604
rect 2724 2570 2762 2604
rect 2796 2570 2834 2604
rect 2868 2570 2906 2604
rect 2940 2570 2978 2604
rect 3012 2570 3050 2604
rect 3084 2570 3122 2604
rect 3156 2570 3194 2604
rect 3228 2570 3266 2604
rect 3300 2570 3338 2604
rect 3372 2570 3410 2604
rect 3444 2570 3482 2604
rect 3516 2570 3554 2604
rect 3588 2570 3626 2604
rect 3660 2570 3698 2604
rect 3732 2598 7740 2604
rect 7774 2598 7812 2632
rect 7846 2598 7884 2632
rect 7918 2598 7956 2632
rect 7990 2598 8028 2632
rect 8062 2598 8100 2632
rect 8134 2598 8172 2632
rect 8206 2598 8244 2632
rect 8278 2598 8316 2632
rect 8350 2598 8388 2632
rect 8422 2598 8460 2632
rect 8494 2598 8532 2632
rect 8566 2598 8604 2632
rect 8638 2598 8676 2632
rect 8710 2598 8748 2632
rect 8782 2598 8820 2632
rect 8854 2598 8892 2632
rect 8926 2598 8964 2632
rect 8998 2598 9036 2632
rect 9070 2598 9108 2632
rect 9142 2598 9245 2632
rect 3732 2576 9245 2598
rect 3732 2570 5030 2576
rect -5114 2542 5030 2570
rect 5064 2542 5102 2576
rect 5136 2542 5174 2576
rect 5208 2542 5246 2576
rect 5280 2542 5318 2576
rect 5352 2542 5390 2576
rect 5424 2542 5462 2576
rect 5496 2542 5534 2576
rect 5568 2542 5606 2576
rect 5640 2542 5678 2576
rect 5712 2542 5750 2576
rect 5784 2542 5822 2576
rect 5856 2542 5894 2576
rect 5928 2542 5966 2576
rect 6000 2542 6038 2576
rect 6072 2542 6110 2576
rect 6144 2542 6182 2576
rect 6216 2542 6254 2576
rect 6288 2542 6326 2576
rect 6360 2542 6398 2576
rect 6432 2542 9245 2576
rect -5114 2462 9245 2542
<< via1 >>
rect -4794 5082 -4734 5142
rect -3688 5088 -3628 5148
rect -4730 4882 -4674 5032
rect -4824 2848 -4764 2902
rect -3692 2844 -3632 2898
<< metal2 >>
rect -4794 5148 -4734 5152
rect -3688 5148 -3628 5158
rect -4802 5142 -3688 5148
rect -4802 5090 -4794 5142
rect -4734 5090 -3688 5142
rect -4794 5072 -4734 5082
rect -4696 5042 -4658 5090
rect -3688 5078 -3628 5088
rect -4730 5032 -4658 5042
rect -4674 4884 -4658 5032
rect -4730 4872 -4674 4882
rect -4824 2910 -4764 2912
rect -4836 2902 -3632 2910
rect -4836 2848 -4824 2902
rect -4764 2898 -3632 2902
rect -4764 2848 -3692 2898
rect -4824 2838 -4764 2848
rect -3692 2834 -3632 2844
use sky130_fd_pr__nfet_01v8_ZE46K8  sky130_fd_pr__nfet_01v8_ZE46K8_0
timestamp 1608322001
transform -1 0 -3669 0 -1 3045
box -211 -319 211 319
use via_li_m1  via_li_m1_1
array 0 19 72 0 0 74
timestamp 1607692587
transform 1 0 -4942 0 1 2536
box 4 0 76 74
use via_li_m1  via_li_m1_0
array 0 19 72 0 0 74
timestamp 1607692587
transform 1 0 -4942 0 1 2636
box 4 0 76 74
use sky130_fd_pr__nfet_01v8_YK3456  sky130_fd_pr__nfet_01v8_YK3456_0
timestamp 1608249442
transform -1 0 -4795 0 -1 3024
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_9TXQ83  sky130_fd_pr__nfet_01v8_9TXQ83_1
timestamp 1608229483
transform 1 0 9023 0 1 3574
box -211 -264 211 264
use sky130_fd_pr__nfet_01v8_R7545W  sky130_fd_pr__nfet_01v8_R7545W_0
timestamp 1608229183
transform 1 0 8231 0 1 3560
box -211 -330 211 330
use via_li_m1  via_li_m1_4
array 0 13 72 0 0 74
timestamp 1607692587
transform 1 0 8148 0 1 3136
box 4 0 76 74
use inverter  inverter_1
array 0 20 569 0 0 858
timestamp 1608329555
transform 1 0 990 0 1 3228
box -5393 252 -4418 1124
use sky130_fd_pr__pfet_01v8_373K6R  sky130_fd_pr__pfet_01v8_373K6R_0
timestamp 1608255150
transform 1 0 9023 0 1 4269
box -211 -327 211 327
use sky130_fd_pr__pfet_01v8_3FZUWK  sky130_fd_pr__pfet_01v8_3FZUWK_0
timestamp 1608254796
transform 1 0 8231 0 1 4426
box -211 -436 211 459
use sky130_fd_pr__pfet_01v8_35M7SK  sky130_fd_pr__pfet_01v8_35M7SK_0
timestamp 1608326616
transform -1 0 -4765 0 1 4961
box -211 -128 211 188
use sky130_fd_pr__pfet_01v8_3D5K6R  sky130_fd_pr__pfet_01v8_3D5K6R_0
timestamp 1608253231
transform 1 0 -3667 0 1 4954
box -211 -324 211 324
use via_li_m1  via_li_m1_3
array 0 19 72 0 0 74
timestamp 1607692587
transform 1 0 -4914 0 1 5286
box 4 0 76 74
use via_li_m1  via_li_m1_2
array 0 19 72 0 0 74
timestamp 1607692587
transform 1 0 -4906 0 1 5386
box 4 0 76 74
<< labels >>
rlabel metal1 9050 3886 9347 3920 1 out_vco
rlabel metal1 8258 3886 8689 3922 1 out_ring
rlabel metal1 -5114 2462 -3040 2804 1 vss
rlabel metal1 -5122 5198 -2718 5516 1 vdd
rlabel metal2 -4764 2848 -3692 2910 1 in
rlabel space -4324 3520 8202 3624 1 9
rlabel metal1 -4314 4172 7952 4352 1 10
rlabel metal2 -4734 5090 -3688 5148 1 5
<< end >>
